module ss_core (

);



endmodule