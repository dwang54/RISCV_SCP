module top (

);



endmodule