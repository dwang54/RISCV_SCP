module SS_Core (

);



endmodule